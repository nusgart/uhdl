// <MODULE> --- <SHORT DESCRIPTION>
//
// <LONG DESCRIPTION>
//
// <FOR ORIGINAL FILES THAT ARE BASED ON ORIGINAL CADR SCHEMATICS:>
// HISTORY:
//
//   (20YY-MM-DD HH:mm:ss AUTHOR) COMMENT

`timescale 1ns/1ps
`default_nettype none

module <MODULE>(/*AUTOARG*/);

   // Inputs and outputs.

   /*AUTOINPUT*/
   /*AUTOOUTPUT*/
   /*AUTOINOUT*/

   ////////////////////////////////////////////////////////////////////////////////

   /*AUTOREG*/
   /*AUTOWIRE*/
   // Add extra wires and registers here, in lexiographical order.

   ////////////////////////////////////////////////////////////////////////////////

   /// Start writing here.

endmodule

`default_nettype wire

// Local Variables:
// verilog-library-directories: ("..")
// End:
