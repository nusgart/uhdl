// cadr.vh --- global definitions
