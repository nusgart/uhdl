// CLOCK1 --- MASTER CLOCK
//
// ---!!! Remove this module.
//
// History:
//
//   (1978-08-30 20:55:32 TK) Initial.

`timescale 1ns/1ps
`default_nettype none

module CLOCK1
  ();

endmodule

`default_nettype wire

// Local Variables:
// verilog-library-directories: ("../..")
// End:
