// BCTERM --- BUSINT CABLE TERMINATION
//
// ---!!! Remove this module.
//
// History:
//
//   (1978-06-21 02:30:59) Initial.

`timescale 1ns/1ps
`default_nettype none

module BCTERM
  ();

endmodule

`default_nettype wire

// Local Variables:
// verilog-library-directories: ("..")
// End:
