module SPCLCH (spc, spco);

   output [18:0] spc;
   input [18:0]  spco;

   // mux SPC
   assign spc = spco;

endmodule
