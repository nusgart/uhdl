// CLOCK2 --- MASTER CLOCK
//
// ---!!! Remove this module.
//
// History:
//
//   (1978-10-11 15:34:47 TK) Initial.

`timescale 1ns/1ps
`default_nettype none

module CLOCK2(/*AUTOARG*/);

endmodule

`default_nettype wire

// Local Variables:
// verilog-library-directories: ("../..")
// End:
