// CPINS --- BUS INTERFACE CABLES
//
// ---!!! Remove this module.
//
// History:
//
//   (1978-08-22 11:23:08 TK) Initial.

`timescale 1ns/1ps
`default_nettype none

module CPINS
  ();

endmodule

`default_nettype wire

// Local Variables:
// verilog-library-directories: ("..")
// End:
