// part_32x32prom_maskright.v --- 32x32 ROM
//
// Used by MSKG4 (RIGHT).

module part_32x32prom_maskright(clk, addr, q);

   input clk;
   input [4:0] addr;
   output [31:0] q;

   ////////////////////////////////////////////////////////////////////////////////

   reg [31:0] q;

   ////////////////////////////////////////////////////////////////////////////////

   always @(posedge clk)
     case (addr)
       5'o00: q = 32'b11111111111111111111111111111111;
       5'o01: q = 32'b11111111111111111111111111111110;
       5'o02: q = 32'b11111111111111111111111111111100;
       5'o03: q = 32'b11111111111111111111111111111000;
       5'o04: q = 32'b11111111111111111111111111110000;
       5'o05: q = 32'b11111111111111111111111111100000;
       5'o06: q = 32'b11111111111111111111111111000000;
       5'o07: q = 32'b11111111111111111111111110000000;
       5'o10: q = 32'b11111111111111111111111100000000;
       5'o11: q = 32'b11111111111111111111111000000000;
       5'o12: q = 32'b11111111111111111111110000000000;
       5'o13: q = 32'b11111111111111111111100000000000;
       5'o14: q = 32'b11111111111111111111000000000000;
       5'o15: q = 32'b11111111111111111110000000000000;
       5'o16: q = 32'b11111111111111111100000000000000;
       5'o17: q = 32'b11111111111111111000000000000000;
       5'o20: q = 32'b11111111111111110000000000000000;
       5'o21: q = 32'b11111111111111100000000000000000;
       5'o22: q = 32'b11111111111111000000000000000000;
       5'o23: q = 32'b11111111111110000000000000000000;
       5'o24: q = 32'b11111111111100000000000000000000;
       5'o25: q = 32'b11111111111000000000000000000000;
       5'o26: q = 32'b11111111110000000000000000000000;
       5'o27: q = 32'b11111111100000000000000000000000;
       5'o30: q = 32'b11111111000000000000000000000000;
       5'o31: q = 32'b11111110000000000000000000000000;
       5'o32: q = 32'b11111100000000000000000000000000;
       5'o33: q = 32'b11111000000000000000000000000000;
       5'o34: q = 32'b11110000000000000000000000000000;
       5'o35: q = 32'b11100000000000000000000000000000;
       5'o36: q = 32'b11000000000000000000000000000000;
       5'o37: q = 32'b10000000000000000000000000000000;
     endcase

endmodule
