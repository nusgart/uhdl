// CAPS --- BYPASS CAPACITORS
//
// ---!!! Remove this module.
//
// History:
//
//   (1978-02-16 04:36:34 TK) Initial.

`timescale 1ns/1ps
`default_nettype none

module CAPS
  ();

endmodule

`default_nettype wire

// Local Variables:
// verilog-library-directories: ("..")
// End:
