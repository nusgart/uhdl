// SPY2 --- PDP11 EXAMINE (A, M, FLAG2)
//
// ---!!! Add description.
//
// History:
//
//   (20YY-MM-DD HH:mm:ss BRAD) Converted to Verilog; merge of ???
//	and ???.
//	???: Nets added.
//	???: Nets removed.
//   (1978-08-16 05:46:29 TK) Initial.

`timescale 1ns/1ps
`default_nettype none

module SPY2(/*AUTOARG*/);

endmodule

`default_nettype wire

// Local Variables:
// verilog-library-directories: ("..")
// End:
