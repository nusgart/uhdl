// IOR
//
// TK		CADR	INST. MODIFY OR

module IOR(iob, i, ob);

   input [31:0] ob;
   input [48:0] i;
   output [47:0] iob;

   ////////////////////////////////////////////////////////////////////////////////

   // iob 47 46 45 44 43 42 41 40 39 38 37 36 35 34 33 32 31 30 29 28 27 26
   // i   47 46 45 44 43 42 41 40 39 38 37 36 35 34 33 32 31 30 29 28 27 26
   // ob  21 20 19 18 17 16 15 14 13 12 11 10 9  8  7  6  5  4  3  2  1  0

   // iob 25 24 ... 1  0
   // i   25 24 ... 1  0
   // ob  25 24 ... 1  0

   assign iob = i[47:0] | { ob[21:0], ob[25:0] };

endmodule
