// MBCPIN --- BUS INTERFACE CABLES
//
// ---!!! Remove this module.
//
// History:
//
//   (1978-08-16 09:01:25 TK) Initial.

`timescale 1ns/1ps
`default_nettype none

module MBCPIN
  ();

endmodule

`default_nettype wire

// Local Variables:
// verilog-library-directories: ("../..")
// End:
