// ICAPS --- BYPASS CAPACITORS
//
// ---!!! Remove this module.
//
// History:
//
//   (1978-10-11 15:21:38 TK) Initial.

`timescale 1ns/1ps
`default_nettype none

module ICAPS
  ();

endmodule

`default_nettype wire

// Local Variables:
// verilog-library-directories: ("../..")
// End:
