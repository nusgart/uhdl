// IWRPAR --- IWR PARITY
//
// ---!!! Remove this module; we don't need parity.
//
// History:
//
//   (1978-01-26 22:54:41 TK) Initial.

`timescale 1ns/1ps
`default_nettype none

module IWRPAR
  ();

endmodule

`default_nettype wire

// Local Variables:
// verilog-library-directories: ("../..")
// End:
