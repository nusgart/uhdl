// SPY4 --- PDP11 EXAMINE (OPC, FLAG1, PC)
//
// ---!!! Add description.
//
// History:
//
//   (20YY-MM-DD HH:mm:ss BRAD) Converted to Verilog; merge of ???
//	and ???.
//	???: Nets added.
//	???: Nets removed.
//   (1978-08-16 09:04:42 TK) Initial.

`timescale 1ns/1ps
`default_nettype none

module SPY4(/*AUTOARG*/);

endmodule

`default_nettype wire

// Local Variables:
// verilog-library-directories: ("../..")
// End:
