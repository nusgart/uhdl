// SPY1 --- PDP11 EXAMINE (IR, OB)
//
// ---!!! Add description.
//
// History:
//
//   (20YY-MM-DD HH:mm:ss BRAD) Converted to Verilog; merge of ???
//	and ???.
//	???: Nets added.
//	???: Nets removed.
//   (1978-01-24 13:43:13 TK) Initial.

`timescale 1ns/1ps
`default_nettype none

module SPY1
  ();

endmodule

`default_nettype wire

// Local Variables:
// verilog-library-directories: ("..")
// End:
