// STAT --- STATISTICS COUNTER
//
// ---!!! Add description.
//
// History:
//
//   (20YY-MM-DD HH:mm:ss BRAD) Converted to Verilog.
//	???: Nets added.
//	???: Nets removed.
//   (1978-06-24 04:25:26 TK) Initial.

`timescale 1ns/1ps
`default_nettype none

module STAT
  ();

endmodule

`default_nettype wire

// Local Variables:
// verilog-library-directories: ("../../..")
// End:
