 `define ISE

`define x512Mb
`define FULL_MEM
`define sg5
`define x16

`define use_ucode_ram

