// CLOCKD --- CLOCK DISTRIBUTION
//
// ---!!! Remove this module.
//
// History:
//
//   (1978-05-08 07:04:53 TK) Initial.

`timescale 1ns/1ps
`default_nettype none

module CLOCKD(/*AUTOARG*/);

endmodule

`default_nettype wire

// Local Variables:
// verilog-library-directories: ("..")
// End:
