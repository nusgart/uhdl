// APAR --- A&M PARITY
//
// ---!!! Remove this module.
//
// History:
//
//   (1978-01-23 10:40:10 TK) Initial.

`timescale 1ns/1ps
`default_nettype none

module APAR(/*AUTOARG*/);

endmodule

`default_nettype wire

// Local Variables:
// verilog-library-directories: ("..")
// End:
