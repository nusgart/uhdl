// SPCPAR --- SPC MEMORY PARITY
//
// ---!!! Remove this module; we don't need parity.
//
// History:
//
//   (1978-01-23 06:33:37 TK) Initial.

`timescale 1ns/1ps
`default_nettype none

module SPCPAR
  ();

endmodule

`default_nettype wire

// Local Variables:
// verilog-library-directories: ("..")
// End:
