// IPAR --- IR PARITY
//
// ---!!! Remove this module; we don't need parity.
//
// History:
//
//   (1978-01-22 12:22:55 TK) Initial.

`timescale 1ns/1ps
`default_nettype none

module IPAR
  ();

endmodule

`default_nettype wire

// Local Variables:
// verilog-library-directories: ("..")
// End:
