// BCPINS --- BUS INTERFACE CABLES
//
// ---!!! Remove this module.
//
// History:
//
//   (1978-08-16 05:02:33 TK) Initial.

`timescale 1ns/1ps
`default_nettype none

module BCPINS(/*AUTOARG*/);

endmodule

`default_nettype wire

// Local Variables:
// verilog-library-directories: ("..")
// End:
