// cadr.vh --- global definitions
`define enable_vga
`define enable_ps2
`define enable_mmc
`define enable_spy_port
`define ISE