// MCPINS --- CONNECTOR PINS
//
// ---!!! Remove this module.
//
// History:
//
//   (1978-08-22 11:29:58 TK) Initial.

`timescale 1ns/1ps
`default_nettype none

module MCPINS
  ();

endmodule

`default_nettype wire

// Local Variables:
// verilog-library-directories: ("../..")
// End:
